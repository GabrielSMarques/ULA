-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

library ieee;
use ieee.std_logic_1164.all;
library altera;
use altera.altera_syn_attributes.all;

entity sdProjectPinPlaner2 is
	port
	(
		A0 : in std_logic;
		A1 : in std_logic;
		A2 : in std_logic;
		A3 : in std_logic;
		A4 : in std_logic;
		ADEZA : out std_logic;
		ADEZB : out std_logic;
		ADEZC : out std_logic;
		ADEZD : out std_logic;
		ADEZE : out std_logic;
		ADEZF : out std_logic;
		ADEZG : out std_logic;
		ASIGNAL : out std_logic;
		AUNIA : out std_logic;
		AUNIB : out std_logic;
		AUNIC : out std_logic;
		AUNID : out std_logic;
		AUNIE : out std_logic;
		AUNIF : out std_logic;
		AUNIG : out std_logic;
		B0 : in std_logic;
		B1 : in std_logic;
		B2 : in std_logic;
		B3 : in std_logic;
		B4 : in std_logic;
		BDEZA : out std_logic;
		BDEZB : out std_logic;
		BDEZC : out std_logic;
		BDEZD : out std_logic;
		BDEZE : out std_logic;
		BDEZF : out std_logic;
		BDEZG : out std_logic;
		BSIGNAL : out std_logic;
		BUNIA : out std_logic;
		BUNIB : out std_logic;
		BUNIC : out std_logic;
		BUNID : out std_logic;
		BUNIE : out std_logic;
		BUNIF : out std_logic;
		BUNIG : out std_logic;
		OUTCOMP : out std_logic;
		R0 : out std_logic;
		R1 : out std_logic;
		R2 : out std_logic;
		R3 : out std_logic;
		R4 : out std_logic;
		S0 : in std_logic;
		S1 : in std_logic;
		S2 : in std_logic;
		SIGNAL : out std_logic
	);

end sdProjectPinPlaner2;

architecture ppl_type of sdProjectPinPlaner2 is

begin

end;
